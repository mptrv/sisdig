.title Tensão de Saída em Função da Resistência do LDR

.include "/home/mpt/Documentos/Projetos/kicad-libraries/kicad-spice-library/Models/uncategorized/spice_complete/NATBJT.LIB"
.include "/home/mpt/Documentos/Projetos/sisdig/1.3-laboratorio/projetos/sensor-e-atuador-com-ajuste-digital-de-set-point/simulacoes/mais-didatico/vres.lib"

.save all
.probe alli

.param Vf = 11.3V
.param tb = 10m
.param ts = 5us
.param td = 'ts'

.param Ka=0
.param Kb=0
.param Kc=1
.param Kd=1

.param Va='Vf*Ka'
.param Vb='Vf*Kb'
.param Vc='Vf*Kc'
.param Vd='Vf*Kd'

V1 VCC 0 Vf

VA1 /Ar 0 DC Va AC 0
VB1 /Br 0 DC Vb AC 0
VC1 /Cr 0 DC Vc AC 0
VD1 /Dr 0 DC Vd AC 0

R10 /V+ /Ar 22k
R1 Net-_R1-Pad1_ 0 22k
R2 Net-_R1-Pad1_ /Dr 22k
R4 Net-_R3-Pad1_ /Cr 22k
R8 Net-_R5-Pad1_ /Br 22k
R9 /V+ Net-_R5-Pad1_ 11k
R16 0 /Vsensor 1Meg
XU1 /Vldr /Vsensor VCC 0 /Vsensor LM324N
XU2 /V+ /Vu2- VCC 0 /Vref LM324N
R12 Net-_R12-Pad1_ /Vu2- 100k
R17 /Vu2- 0 270k
R20 /Vcomp /Vs 100k
R19 /Vref /Vcomp 15k
XU3 /Vcomp /Vsensor VCC 0 /Vs LM324N
R21 0 /Vs 1Meg
R5 Net-_R5-Pad1_ Net-_R3-Pad1_ 11k
R3 Net-_R3-Pad1_ Net-_R1-Pad1_ 11k
R6 0 Net-_R11-Pad1_ 4.7k

RP1 Net-_R11-Pad1_ /Vldr 14k
RP2 /Vref Net-_R12-Pad1_ 50k

Rldr /Vldr VCC 10k

.control

	set color2=blue
	set color3=orange
	set color4=green3
	set color5=red
	set xbrushwidth=3

	let ind = 0
	let nimg = 1
	let npontos = 150
	let passo = $&npontos / $&nimg
	
	*** Rldr crescente
	dc Rldr 1k 150k 1k

	*** Rldr decrescente
	dc Rldr 150k 1k -1k


	*** Gráficos Rldr decrescente

	let ind = 150
	setplot dc2

	repeat $&nimg

		plot "/Vref"  "/Vs" "/Vsensor" "/Vcomp" xlabel 'Rldr decrescente (clareando)' xlimit 0 150k ylimit -0.1 12 xindices 1 $&ind

		let ind = ind - $&passo
	
	end

	*** Gráficos Rldr crescente

	let ind = 150
	setplot dc1

	repeat $&nimg

		plot "/Vref"  "/Vs" "/Vsensor" "/Vcomp" xlabel 'Rldr crescente (escurecendo)' xlimit 0 150k ylimit -0.1 12 xindices 1 $&ind

		let ind = ind - $&passo

	end

	*** Gráfico Combinado

	set color2=red
	set color3=orange
	set color4=red
	set color5=orange
	set color6=green3
	set color7=blue

	plot "dc2./VComp" "dc2./Vs" "dc1./Vcomp" "dc1./Vs" "dc1./Vsensor" "dc1./Vref" xlabel 'Rldr crescente e decrescente' xlimit 0 150k ylimit -0.1 12 xindices 1 $&ind


	* (Para listar ids das janelas: wmctrl -l | grep -e "0x.*N/A$")
		  shell wmctrl -i -r "0x04000011" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000024" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000035" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000046" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000057" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000068" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000079" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x0400008a" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x0400009b" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040000ac" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040000bd" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040000ce" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040000df" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040000f0" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000101" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000112" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000123" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000134" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000145" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000156" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000167" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000178" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000189" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x0400019a" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040001ab" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040001bc" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040001cd" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040001de" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040001ef" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000200" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000211" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000222" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000233" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000244" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000255" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000266" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000277" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000288" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000299" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040002aa" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040002bb" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040002cc" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040002dd" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040002ee" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040002ff" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000310" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000321" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000332" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000343" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000354" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000365" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000376" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000387" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x04000398" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040003a9" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040003ba" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040003cb" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040003dc" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040003ed" -e "0,50,50,935,845"
		  shell wmctrl -i -r "0x040003fe" -e "0,50,50,935,845"

.endc

.end
